(* blackbox *) module RAM128(CLK, EN0, VGND, VPWR, A0, Di0, Do0, WE0);
input CLK, EN0, VGND, VPWR;
input [6:0] A0; input [31:0] Di0; input [3:0] WE0; output [31:0] Do0;
endmodule
(* blackbox *) module RAM256(VPWR, VGND, CLK, WE0, EN0, A0, Di0, Do0);
inout VPWR, VGND; input CLK, EN0;
input [7:0] A0; input [31:0] Di0; input [3:0] WE0; output [31:0] Do0;
endmodule
(* blackbox *) module dummy_por(vdd3v3, vdd1v8, vss3v3, vss1v8, porb_h, porb_l, por_l);
inout vdd3v3, vdd1v8, vss3v3, vss1v8;
output porb_h, porb_l, por_l;
endmodule
